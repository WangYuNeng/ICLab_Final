`ifndef _ECCDefine_VH_
`define _ECCDefine_VH_

`define MAX_BITS 256
`define MAX_REG  7  // lg(MAX_BITS) - 1

// operating mode
`define BITS256 2'b11
`define BITS128 2'b10
`define BITS64  2'b01
`define BITS32  2'b00

`endif