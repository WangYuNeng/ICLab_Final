`ifndef _ECCDefine_VH_
`define _ECCDefine_VH_

`define MAX_BITS 130
`define MAX_REG  6  // lg(MAX_BITS) - 1

// operating mode
`define BITS128 2'b11
`define BITS64  2'b10
`define BITS32  2'b01
`define BITS16  2'b00

`endif
